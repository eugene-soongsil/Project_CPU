module ExcuteRegister(
    input           clk, reset, enalbe,
    input   [11:0]  
    output
    
);


endmodule