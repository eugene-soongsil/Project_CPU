module Team4_CPU(
    input               clk, reset,
    output  [15:0]      DataOut
);




endmodule