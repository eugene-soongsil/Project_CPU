module Team4_CPU(
    input   i_clk,
    input   i_reset,
    input   i_stop,
    output  [3:0]o_write_add,
    output  [7:0]o_write_data
);




endmodule