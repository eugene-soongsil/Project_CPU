module ProgramCounter(
    input           i_clk,
    input           i_reset,
    input           enable,
    input  [11:0]   i_pcOld
    output [11:0]   o_pcNew,
);

reg     [11:0]      r_pcNew;

always@(posedge i_clk or negedge i_reset)begin
    if(~i_reset)
        r_pcNew <= 0;
    else if(~enable)
        r_pcNew <= i_pcOld;
end

assign o_pcNew = r_pcNew;

endmodule