module ControlUnit(
    input [3:0] i_opcode,
    input       i_reset,
    output      o_stallF,
    output      o_stallD,
    output      o_stallE,
    output      o_write_en,
    output      o_setPC,
    output      
);



endmodule