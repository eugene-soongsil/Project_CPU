module DataPath(

);


endmodule